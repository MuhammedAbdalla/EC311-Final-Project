// Display text on the 7-segment display.
// a series of encoded letters to display onto the seven_segments
module text_display();

endmodule