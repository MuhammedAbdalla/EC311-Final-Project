// Aryaman and Aya


module rand_num_generator();

endmodule