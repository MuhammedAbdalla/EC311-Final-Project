// TOP LEVEL MODULE
// INSTANTIATES ALL MODULES

module top(clk, reset);


endmodule