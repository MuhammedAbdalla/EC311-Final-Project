// Track the points via a counter. Decimal output

module points();

endmodule
