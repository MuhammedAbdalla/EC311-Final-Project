// Utilized the rand_num_generator to light up the LED correspondin 
// to integer value 0 <= I <= 15


module choose_mole();

endmodule  